
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MIPSCPU is
  port(clk:in std_logic; Overflow:out std_logic);
end MIPSCPU;

--This is where all the port mapping jawns are
  
  
  architecture Behavorial of MIPSCPU is
  begin
    
  
  end Behavorial;